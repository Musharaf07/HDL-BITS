// Note the Verilog-1995 module declaration syntax here:
module top_module(clk, reset, in, out);
    input clk;
    input reset;    // Synchronous reset to state B
    input in;
    output out;//  
    reg out;

    parameter A = 0, B = 1;
    reg present_state, next_state;

    always @(posedge clk) begin
        if (reset) begin 
            present_state <= B;
        end
        else
            present_state <= next_state;
        end
        
        always@(*)begin
            case(present_state)
                A : next_state = in ? A : B;
                B : next_state = in ? B : A;
                default next_state = A ;
            endcase 
        end
        assign out = (present_state==B);
        endmodule
