module top_module ( input a, input b, output out );
  
    mod_a instance0 (a,b,out);

endmodule
